module bin_to_bcd_14 (
    input[13:0] b, //���14'b11_1111_1111_1111=16383��9999=14'b10_0111_0000_1111
    output reg[16:0] p //16383��ӦBCD����17λ��9999��ӦBCD��Ϊ16'b1001_1001_1001_1001 
);
    //��4��3����ԭ��û��
    reg[32:0] z; //����Ϊɶ33λ
    integer i;

    always@(*) begin
        for(i=0;i<=32;i=i+1) z[i]=0;    
        z[16:3]=b; //ֱ�Ӱ�b����3λ��
        repeat(11) //һ��14�Σ�ǰ���Ѿ��ƶ���3��
        begin
            if(z[17:14]>4) //�����λ����4
                z[17:14]=z[17:14]+3;
            else;
            if(z[21:18]>4) //���ʮλ����4
                z[21:18]=z[21:18]+3;
            else;
            if(z[25:22]>4) //�����λ����4
                z[25:22]=z[25:22]+3;
            else;
            if(z[29:26]>4) //���ǧλ����4
                z[29:26]=z[29:26]+3;
            else;
            z[32:1]=z[31:0]; //����һλ
        end
        p=z[30:14]; //���2λû��
    end
    
endmodule