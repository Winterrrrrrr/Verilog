module bin_to_bcd_14 (
    input[13:0] b, //���ֵΪ14'b11_1111_1111_1111=16383�����������ʾ�����ֵΪ9999=14'b10_0111_0000_1111
    output reg[16:0] p //16383��ӦBCD����17λ��9999��ӦBCD��Ϊ16'b1001_1001_1001_1001����14λ 
);
    //��CSDN�ϲ鵽�Ľ�������ת��Ϊ8421���һ�ּȸ�Ч�ֽ�ʡ��Դ�ķ���
    //��������Ϊ��4��3��������ԭ�����ϵĸ��಩�Ͷ����ɲ��꣬�Ҹ��˲��Ǻܶ�
    //ֻ֪���������õ������ĳλ����4����2���Ӧ��8421��ͱ����λ�������ǰ��3��֤����ȷ������λ�ź�
    //�����Ǿ���ʵ�ִ���

    reg[30:0] z; //�������ƴ洢�����14λ��Ȼ��ͨ��ѭ�����ƣ��������17λ����BCD��
    integer i;

    always@(*) begin
        for(i=0;i<=30;i=i+1) z[i]=0;    
        z[16:3]=b; //ֱ�Ӱ�b����3λ��
        repeat(11) //һ��14λ������Ҫ��λ14�Σ�ǰ���Ѿ��ƶ���3�Σ�������������λ11��
        begin
            if(z[17:14]>4) //�����λ����4
                z[17:14]=z[17:14]+3;
            else;
            if(z[21:18]>4) //���ʮλ����4
                z[21:18]=z[21:18]+3;
            else;
            if(z[25:22]>4) //�����λ����4
                z[25:22]=z[25:22]+3;
            else;
            if(z[29:26]>4) //���ǧλ����4
                z[29:26]=z[29:26]+3;
            else;
            z[30:1]=z[29:0]; //����һλ
        end
        p=z[30:14]; 
    end
    
endmodule