module binbcd8 (
    input[7:0] b,
    output reg[9:0] p //8λ�����������1111_1111����Ӧ255��BCD����10 0101 0101
);
    //��4��3����ԭ��û��
    reg[17:0] z;
    always@(*) begin
        z=18'b00_0000_0000_0000_0000;
        z[10:3]=b; //ֱ�Ӱ�b����3λ��
        repeat(5) //һ��8�Σ�ǰ���Ѿ��ƶ���5��
        begin
            if(z[11:8]>4)
                z[11:8]=z[11:8]+3;
            else;
            if(z[15:12]>4)
                z[15:12]=z[15:12]+3;
            else;
            //��ߵ�4λ�϶��������4����Ϊ��255��ֻ��0010
            z[17:1]=z[16:0]; //����һλ
        end
        p=z[17:8];
    end
    
endmodule